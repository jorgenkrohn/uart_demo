library ieee;
use ieee.std_logic_1164.all;

package uart_vvc_tb_pkg is

  constant C_TX_IDX   : natural := 0;
  constant C_RX_IDX   : natural := 1;
  constant C_UART_IDX : natural := 0;
  
end package uart_vvc_tb_pkg;
